
module progmem (
    // Closk & reset
    input wire clk,
    input wire rstn,

    // PicoRV32 bus interface
    input  wire        valid,
    output wire        ready,
    input  wire [31:0] addr,
    output wire [31:0] rdata
);

  // ============================================================================

  localparam MEM_SIZE_BITS = 10;  // In 32-bit words
  localparam MEM_SIZE = 1 << MEM_SIZE_BITS;
  localparam MEM_ADDR_MASK = 32'h0010_0000;

  // ============================================================================

  wire [MEM_SIZE_BITS-1:0] mem_addr;
  reg  [             31:0] mem_data;
  reg  [             31:0] mem      [0:MEM_SIZE];

  initial begin
    mem['h0000] <= 32'h00000093;
    mem['h0001] <= 32'h00000193;
    mem['h0002] <= 32'h00000213;
    mem['h0003] <= 32'h00000293;
    mem['h0004] <= 32'h00000313;
    mem['h0005] <= 32'h00000393;
    mem['h0006] <= 32'h00000413;
    mem['h0007] <= 32'h00000493;
    mem['h0008] <= 32'h00000513;
    mem['h0009] <= 32'h00000593;
    mem['h000A] <= 32'h00000613;
    mem['h000B] <= 32'h00000693;
    mem['h000C] <= 32'h00000713;
    mem['h000D] <= 32'h00000793;
    mem['h000E] <= 32'h00000813;
    mem['h000F] <= 32'h00000893;
    mem['h0010] <= 32'h00000913;
    mem['h0011] <= 32'h00000993;
    mem['h0012] <= 32'h00000A13;
    mem['h0013] <= 32'h00000A93;
    mem['h0014] <= 32'h00000B13;
    mem['h0015] <= 32'h00000B93;
    mem['h0016] <= 32'h00000C13;
    mem['h0017] <= 32'h00000C93;
    mem['h0018] <= 32'h00000D13;
    mem['h0019] <= 32'h00000D93;
    mem['h001A] <= 32'h00000E13;
    mem['h001B] <= 32'h00000E93;
    mem['h001C] <= 32'h00000F13;
    mem['h001D] <= 32'h00000F93;
    mem['h001E] <= 32'h00000513;
    mem['h001F] <= 32'h00000593;
    mem['h0020] <= 32'h00B52023;
    mem['h0021] <= 32'h00450513;
    mem['h0022] <= 32'hFE254CE3;
    mem['h0023] <= 32'h00001517;
    mem['h0024] <= 32'h99C50513;
    mem['h0025] <= 32'h00000593;
    mem['h0026] <= 32'h00000613;
    mem['h0027] <= 32'h00C5DC63;
    mem['h0028] <= 32'h00052683;
    mem['h0029] <= 32'h00D5A023;
    mem['h002A] <= 32'h00450513;
    mem['h002B] <= 32'h00458593;
    mem['h002C] <= 32'hFEC5C8E3;
    mem['h002D] <= 32'h00000513;
    mem['h002E] <= 32'h00000593;
    mem['h002F] <= 32'h00B55863;
    mem['h0030] <= 32'h00052023;
    mem['h0031] <= 32'h00450513;
    mem['h0032] <= 32'hFEB54CE3;
    mem['h0033] <= 32'h008000EF;
    mem['h0034] <= 32'h0000006F;
    mem['h0035] <= 32'hFA010113;
    mem['h0036] <= 32'h04112E23;
    mem['h0037] <= 32'h04812C23;
    mem['h0038] <= 32'h06010413;
    mem['h0039] <= 32'h001017B7;
    mem['h003A] <= 32'hA0478793;
    mem['h003B] <= 32'h0007A603;
    mem['h003C] <= 32'h0047A683;
    mem['h003D] <= 32'h0087A703;
    mem['h003E] <= 32'hFEC42023;
    mem['h003F] <= 32'hFED42223;
    mem['h0040] <= 32'hFEE42423;
    mem['h0041] <= 32'h00C7D783;
    mem['h0042] <= 32'hFEF41623;
    mem['h0043] <= 32'hFA040713;
    mem['h0044] <= 32'hFE040793;
    mem['h0045] <= 32'h00070613;
    mem['h0046] <= 32'h00D00593;
    mem['h0047] <= 32'h00078513;
    mem['h0048] <= 32'h7FC000EF;
    mem['h0049] <= 32'h00000013;
    mem['h004A] <= 32'h05C12083;
    mem['h004B] <= 32'h05812403;
    mem['h004C] <= 32'h06010113;
    mem['h004D] <= 32'h00008067;
    mem['h004E] <= 32'hFE010113;
    mem['h004F] <= 32'h00812E23;
    mem['h0050] <= 32'h02010413;
    mem['h0051] <= 32'h00050793;
    mem['h0052] <= 32'hFEB42423;
    mem['h0053] <= 32'hFEF407A3;
    mem['h0054] <= 32'hFEF44783;
    mem['h0055] <= 32'h0047D793;
    mem['h0056] <= 32'h0FF7F793;
    mem['h0057] <= 32'h00F7F793;
    mem['h0058] <= 32'h00101737;
    mem['h0059] <= 32'hA1470713;
    mem['h005A] <= 32'h00F707B3;
    mem['h005B] <= 32'h0007C703;
    mem['h005C] <= 32'hFE842783;
    mem['h005D] <= 32'h00E78023;
    mem['h005E] <= 32'hFEF44783;
    mem['h005F] <= 32'h00F7F713;
    mem['h0060] <= 32'hFE842783;
    mem['h0061] <= 32'h00178793;
    mem['h0062] <= 32'h001016B7;
    mem['h0063] <= 32'hA1468693;
    mem['h0064] <= 32'h00E68733;
    mem['h0065] <= 32'h00074703;
    mem['h0066] <= 32'h00E78023;
    mem['h0067] <= 32'hFE842783;
    mem['h0068] <= 32'h00278793;
    mem['h0069] <= 32'h00078023;
    mem['h006A] <= 32'h00000013;
    mem['h006B] <= 32'h01C12403;
    mem['h006C] <= 32'h02010113;
    mem['h006D] <= 32'h00008067;
    mem['h006E] <= 32'hF8010113;
    mem['h006F] <= 32'h06812E23;
    mem['h0070] <= 32'h08010413;
    mem['h0071] <= 32'hF8A42623;
    mem['h0072] <= 32'hF8B42423;
    mem['h0073] <= 32'hFE042623;
    mem['h0074] <= 32'hFE042423;
    mem['h0075] <= 32'h0BC0006F;
    mem['h0076] <= 32'hFE842783;
    mem['h0077] <= 32'h00279793;
    mem['h0078] <= 32'hFF078793;
    mem['h0079] <= 32'h008787B3;
    mem['h007A] <= 32'hFA07A223;
    mem['h007B] <= 32'hFE042223;
    mem['h007C] <= 32'h0880006F;
    mem['h007D] <= 32'hFE842783;
    mem['h007E] <= 32'h00279793;
    mem['h007F] <= 32'hFF078793;
    mem['h0080] <= 32'h008787B3;
    mem['h0081] <= 32'hFA47A783;
    mem['h0082] <= 32'h00879713;
    mem['h0083] <= 32'hFE842783;
    mem['h0084] <= 32'h00279793;
    mem['h0085] <= 32'hFF078793;
    mem['h0086] <= 32'h008787B3;
    mem['h0087] <= 32'hFAE7A223;
    mem['h0088] <= 32'hFE842783;
    mem['h0089] <= 32'h00279793;
    mem['h008A] <= 32'hFF078793;
    mem['h008B] <= 32'h008787B3;
    mem['h008C] <= 32'hFA47A783;
    mem['h008D] <= 32'hFE842703;
    mem['h008E] <= 32'h00271693;
    mem['h008F] <= 32'hFE442703;
    mem['h0090] <= 32'h00E68733;
    mem['h0091] <= 32'h00070693;
    mem['h0092] <= 32'hF8842703;
    mem['h0093] <= 32'h00D70733;
    mem['h0094] <= 32'h00074703;
    mem['h0095] <= 32'h00E7E733;
    mem['h0096] <= 32'hFE842783;
    mem['h0097] <= 32'h00279793;
    mem['h0098] <= 32'hFF078793;
    mem['h0099] <= 32'h008787B3;
    mem['h009A] <= 32'hFAE7A223;
    mem['h009B] <= 32'hFE442783;
    mem['h009C] <= 32'h00178793;
    mem['h009D] <= 32'hFEF42223;
    mem['h009E] <= 32'hFE442703;
    mem['h009F] <= 32'h00300793;
    mem['h00A0] <= 32'hF6E7DAE3;
    mem['h00A1] <= 32'hFE842783;
    mem['h00A2] <= 32'h00178793;
    mem['h00A3] <= 32'hFEF42423;
    mem['h00A4] <= 32'hFE842703;
    mem['h00A5] <= 32'h00F00793;
    mem['h00A6] <= 32'hF4E7D0E3;
    mem['h00A7] <= 32'hFEC42783;
    mem['h00A8] <= 32'hFEC42703;
    mem['h00A9] <= 32'h00E7C78B;
    mem['h00AA] <= 32'hFEF42623;
    mem['h00AB] <= 32'hFE042023;
    mem['h00AC] <= 32'h0380006F;
    mem['h00AD] <= 32'hFE042783;
    mem['h00AE] <= 32'h00279793;
    mem['h00AF] <= 32'hFF078793;
    mem['h00B0] <= 32'h008787B3;
    mem['h00B1] <= 32'hFA47A783;
    mem['h00B2] <= 32'hFCF42A23;
    mem['h00B3] <= 32'hFD442783;
    mem['h00B4] <= 32'hFE042703;
    mem['h00B5] <= 32'h00E7878B;
    mem['h00B6] <= 32'hFEF42623;
    mem['h00B7] <= 32'hFE042783;
    mem['h00B8] <= 32'h00178793;
    mem['h00B9] <= 32'hFEF42023;
    mem['h00BA] <= 32'hFE042703;
    mem['h00BB] <= 32'h00F00793;
    mem['h00BC] <= 32'hFCE7D2E3;
    mem['h00BD] <= 32'hF8C42783;
    mem['h00BE] <= 32'h0447A703;
    mem['h00BF] <= 32'h00100793;
    mem['h00C0] <= 32'h00F71C63;
    mem['h00C1] <= 32'hFEC42783;
    mem['h00C2] <= 32'hFEC42703;
    mem['h00C3] <= 32'h00E7978B;
    mem['h00C4] <= 32'hFEF42623;
    mem['h00C5] <= 32'h0140006F;
    mem['h00C6] <= 32'hFEC42783;
    mem['h00C7] <= 32'hFEC42703;
    mem['h00C8] <= 32'h00E7A78B;
    mem['h00C9] <= 32'hFEF42623;
    mem['h00CA] <= 32'hFC042E23;
    mem['h00CB] <= 32'h03C0006F;
    mem['h00CC] <= 32'hFEC42783;
    mem['h00CD] <= 32'hFDC42703;
    mem['h00CE] <= 32'h00E7B78B;
    mem['h00CF] <= 32'hFCF42C23;
    mem['h00D0] <= 32'hF8C42703;
    mem['h00D1] <= 32'hFDC42783;
    mem['h00D2] <= 32'h01478793;
    mem['h00D3] <= 32'h00279793;
    mem['h00D4] <= 32'h00F707B3;
    mem['h00D5] <= 32'hFD842703;
    mem['h00D6] <= 32'h00E7A023;
    mem['h00D7] <= 32'hFDC42783;
    mem['h00D8] <= 32'h00178793;
    mem['h00D9] <= 32'hFCF42E23;
    mem['h00DA] <= 32'hFDC42703;
    mem['h00DB] <= 32'h00700793;
    mem['h00DC] <= 32'hFCE7D0E3;
    mem['h00DD] <= 32'h00000013;
    mem['h00DE] <= 32'h00000013;
    mem['h00DF] <= 32'h07C12403;
    mem['h00E0] <= 32'h08010113;
    mem['h00E1] <= 32'h00008067;
    mem['h00E2] <= 32'hFE010113;
    mem['h00E3] <= 32'h00812E23;
    mem['h00E4] <= 32'h02010413;
    mem['h00E5] <= 32'hFEA42623;
    mem['h00E6] <= 32'hFEC42783;
    mem['h00E7] <= 32'h0407A023;
    mem['h00E8] <= 32'hFEC42783;
    mem['h00E9] <= 32'h0407A223;
    mem['h00EA] <= 32'hFEC42783;
    mem['h00EB] <= 32'h0407A423;
    mem['h00EC] <= 32'hFEC42783;
    mem['h00ED] <= 32'h0407A623;
    mem['h00EE] <= 32'hFEC42783;
    mem['h00EF] <= 32'h0407A823;
    mem['h00F0] <= 32'hFEC42783;
    mem['h00F1] <= 32'h0407AA23;
    mem['h00F2] <= 32'hFEC42783;
    mem['h00F3] <= 32'h0407AC23;
    mem['h00F4] <= 32'hFEC42783;
    mem['h00F5] <= 32'h0407AE23;
    mem['h00F6] <= 32'hFEC42783;
    mem['h00F7] <= 32'h0607A023;
    mem['h00F8] <= 32'hFEC42783;
    mem['h00F9] <= 32'h0607A223;
    mem['h00FA] <= 32'hFEC42783;
    mem['h00FB] <= 32'h0607A423;
    mem['h00FC] <= 32'hFEC42783;
    mem['h00FD] <= 32'h0607A623;
    mem['h00FE] <= 32'h00000013;
    mem['h00FF] <= 32'h01C12403;
    mem['h0100] <= 32'h02010113;
    mem['h0101] <= 32'h00008067;
    mem['h0102] <= 32'hFD010113;
    mem['h0103] <= 32'h02112623;
    mem['h0104] <= 32'h02812423;
    mem['h0105] <= 32'h03010413;
    mem['h0106] <= 32'hFCA42E23;
    mem['h0107] <= 32'hFCB42C23;
    mem['h0108] <= 32'hFCC42A23;
    mem['h0109] <= 32'hFE042623;
    mem['h010A] <= 32'h0BC0006F;
    mem['h010B] <= 32'hFEC42783;
    mem['h010C] <= 32'hFD842703;
    mem['h010D] <= 32'h00F70733;
    mem['h010E] <= 32'hFDC42783;
    mem['h010F] <= 32'h0407A783;
    mem['h0110] <= 32'h00074703;
    mem['h0111] <= 32'hFDC42683;
    mem['h0112] <= 32'h00F687B3;
    mem['h0113] <= 32'h00E78023;
    mem['h0114] <= 32'hFDC42783;
    mem['h0115] <= 32'h0407A783;
    mem['h0116] <= 32'h00178713;
    mem['h0117] <= 32'hFDC42783;
    mem['h0118] <= 32'h04E7A023;
    mem['h0119] <= 32'hFDC42783;
    mem['h011A] <= 32'h0407A703;
    mem['h011B] <= 32'h04000793;
    mem['h011C] <= 32'h06F71463;
    mem['h011D] <= 32'hFDC42783;
    mem['h011E] <= 32'h0447A783;
    mem['h011F] <= 32'h00178713;
    mem['h0120] <= 32'hFDC42783;
    mem['h0121] <= 32'h04E7A223;
    mem['h0122] <= 32'hFDC42783;
    mem['h0123] <= 32'h00078593;
    mem['h0124] <= 32'hFDC42503;
    mem['h0125] <= 32'hD25FF0EF;
    mem['h0126] <= 32'hFDC42783;
    mem['h0127] <= 32'h0487A703;
    mem['h0128] <= 32'hDFF00793;
    mem['h0129] <= 32'h00E7FC63;
    mem['h012A] <= 32'hFDC42783;
    mem['h012B] <= 32'h04C7A783;
    mem['h012C] <= 32'h00178713;
    mem['h012D] <= 32'hFDC42783;
    mem['h012E] <= 32'h04E7A623;
    mem['h012F] <= 32'hFDC42783;
    mem['h0130] <= 32'h0487A783;
    mem['h0131] <= 32'h20078713;
    mem['h0132] <= 32'hFDC42783;
    mem['h0133] <= 32'h04E7A423;
    mem['h0134] <= 32'hFDC42783;
    mem['h0135] <= 32'h0407A023;
    mem['h0136] <= 32'hFEC42783;
    mem['h0137] <= 32'h00178793;
    mem['h0138] <= 32'hFEF42623;
    mem['h0139] <= 32'hFEC42783;
    mem['h013A] <= 32'hFD442703;
    mem['h013B] <= 32'hF4E7E0E3;
    mem['h013C] <= 32'h00000013;
    mem['h013D] <= 32'h00000013;
    mem['h013E] <= 32'h02C12083;
    mem['h013F] <= 32'h02812403;
    mem['h0140] <= 32'h03010113;
    mem['h0141] <= 32'h00008067;
    mem['h0142] <= 32'hFD010113;
    mem['h0143] <= 32'h02112623;
    mem['h0144] <= 32'h02812423;
    mem['h0145] <= 32'h03010413;
    mem['h0146] <= 32'hFCA42E23;
    mem['h0147] <= 32'hFCB42C23;
    mem['h0148] <= 32'hFDC42783;
    mem['h0149] <= 32'h0407A783;
    mem['h014A] <= 32'hFEF42623;
    mem['h014B] <= 32'hFDC42783;
    mem['h014C] <= 32'h0407A703;
    mem['h014D] <= 32'h03700793;
    mem['h014E] <= 32'h04E7E663;
    mem['h014F] <= 32'hFEC42783;
    mem['h0150] <= 32'h00178713;
    mem['h0151] <= 32'hFEE42623;
    mem['h0152] <= 32'hFDC42703;
    mem['h0153] <= 32'h00F707B3;
    mem['h0154] <= 32'hF8000713;
    mem['h0155] <= 32'h00E78023;
    mem['h0156] <= 32'h01C0006F;
    mem['h0157] <= 32'hFEC42783;
    mem['h0158] <= 32'h00178713;
    mem['h0159] <= 32'hFEE42623;
    mem['h015A] <= 32'hFDC42703;
    mem['h015B] <= 32'h00F707B3;
    mem['h015C] <= 32'h00078023;
    mem['h015D] <= 32'hFEC42703;
    mem['h015E] <= 32'h03700793;
    mem['h015F] <= 32'hFEE7D0E3;
    mem['h0160] <= 32'h09C0006F;
    mem['h0161] <= 32'hFEC42783;
    mem['h0162] <= 32'h00178713;
    mem['h0163] <= 32'hFEE42623;
    mem['h0164] <= 32'hFDC42703;
    mem['h0165] <= 32'h00F707B3;
    mem['h0166] <= 32'hF8000713;
    mem['h0167] <= 32'h00E78023;
    mem['h0168] <= 32'h01C0006F;
    mem['h0169] <= 32'hFEC42783;
    mem['h016A] <= 32'h00178713;
    mem['h016B] <= 32'hFEE42623;
    mem['h016C] <= 32'hFDC42703;
    mem['h016D] <= 32'h00F707B3;
    mem['h016E] <= 32'h00078023;
    mem['h016F] <= 32'hFEC42703;
    mem['h0170] <= 32'h03F00793;
    mem['h0171] <= 32'hFEE7D0E3;
    mem['h0172] <= 32'hFDC42783;
    mem['h0173] <= 32'h0447A783;
    mem['h0174] <= 32'h00178713;
    mem['h0175] <= 32'hFDC42783;
    mem['h0176] <= 32'h04E7A223;
    mem['h0177] <= 32'hFDC42783;
    mem['h0178] <= 32'h00078593;
    mem['h0179] <= 32'hFDC42503;
    mem['h017A] <= 32'hBD1FF0EF;
    mem['h017B] <= 32'hFE042423;
    mem['h017C] <= 32'h0200006F;
    mem['h017D] <= 32'hFDC42703;
    mem['h017E] <= 32'hFE842783;
    mem['h017F] <= 32'h00F707B3;
    mem['h0180] <= 32'h00078023;
    mem['h0181] <= 32'hFE842783;
    mem['h0182] <= 32'h00178793;
    mem['h0183] <= 32'hFEF42423;
    mem['h0184] <= 32'hFE842703;
    mem['h0185] <= 32'h03700793;
    mem['h0186] <= 32'hFCE7DEE3;
    mem['h0187] <= 32'hFDC42783;
    mem['h0188] <= 32'h0487A703;
    mem['h0189] <= 32'hFDC42783;
    mem['h018A] <= 32'h0407A783;
    mem['h018B] <= 32'h00379793;
    mem['h018C] <= 32'hFFF7C793;
    mem['h018D] <= 32'h00E7FC63;
    mem['h018E] <= 32'hFDC42783;
    mem['h018F] <= 32'h04C7A783;
    mem['h0190] <= 32'h00178713;
    mem['h0191] <= 32'hFDC42783;
    mem['h0192] <= 32'h04E7A623;
    mem['h0193] <= 32'hFDC42783;
    mem['h0194] <= 32'h0487A703;
    mem['h0195] <= 32'hFDC42783;
    mem['h0196] <= 32'h0407A783;
    mem['h0197] <= 32'h00379793;
    mem['h0198] <= 32'h00F70733;
    mem['h0199] <= 32'hFDC42783;
    mem['h019A] <= 32'h04E7A423;
    mem['h019B] <= 32'hFDC42783;
    mem['h019C] <= 32'h0487A783;
    mem['h019D] <= 32'h0FF7F713;
    mem['h019E] <= 32'hFDC42783;
    mem['h019F] <= 32'h02E78FA3;
    mem['h01A0] <= 32'hFDC42783;
    mem['h01A1] <= 32'h0487A783;
    mem['h01A2] <= 32'h0087D793;
    mem['h01A3] <= 32'h0FF7F713;
    mem['h01A4] <= 32'hFDC42783;
    mem['h01A5] <= 32'h02E78F23;
    mem['h01A6] <= 32'hFDC42783;
    mem['h01A7] <= 32'h0487A783;
    mem['h01A8] <= 32'h0107D793;
    mem['h01A9] <= 32'h0FF7F713;
    mem['h01AA] <= 32'hFDC42783;
    mem['h01AB] <= 32'h02E78EA3;
    mem['h01AC] <= 32'hFDC42783;
    mem['h01AD] <= 32'h0487A783;
    mem['h01AE] <= 32'h0187D793;
    mem['h01AF] <= 32'h0FF7F713;
    mem['h01B0] <= 32'hFDC42783;
    mem['h01B1] <= 32'h02E78E23;
    mem['h01B2] <= 32'hFDC42783;
    mem['h01B3] <= 32'h04C7A783;
    mem['h01B4] <= 32'h0FF7F713;
    mem['h01B5] <= 32'hFDC42783;
    mem['h01B6] <= 32'h02E78DA3;
    mem['h01B7] <= 32'hFDC42783;
    mem['h01B8] <= 32'h04C7A783;
    mem['h01B9] <= 32'h0087D793;
    mem['h01BA] <= 32'h0FF7F713;
    mem['h01BB] <= 32'hFDC42783;
    mem['h01BC] <= 32'h02E78D23;
    mem['h01BD] <= 32'hFDC42783;
    mem['h01BE] <= 32'h04C7A783;
    mem['h01BF] <= 32'h0107D793;
    mem['h01C0] <= 32'h0FF7F713;
    mem['h01C1] <= 32'hFDC42783;
    mem['h01C2] <= 32'h02E78CA3;
    mem['h01C3] <= 32'hFDC42783;
    mem['h01C4] <= 32'h04C7A783;
    mem['h01C5] <= 32'h0187D793;
    mem['h01C6] <= 32'h0FF7F713;
    mem['h01C7] <= 32'hFDC42783;
    mem['h01C8] <= 32'h02E78C23;
    mem['h01C9] <= 32'hFDC42783;
    mem['h01CA] <= 32'h0447A783;
    mem['h01CB] <= 32'h00178713;
    mem['h01CC] <= 32'hFDC42783;
    mem['h01CD] <= 32'h04E7A223;
    mem['h01CE] <= 32'hFDC42783;
    mem['h01CF] <= 32'h00078593;
    mem['h01D0] <= 32'hFDC42503;
    mem['h01D1] <= 32'hA75FF0EF;
    mem['h01D2] <= 32'hFE042623;
    mem['h01D3] <= 32'h1AC0006F;
    mem['h01D4] <= 32'hFDC42783;
    mem['h01D5] <= 32'h0507A703;
    mem['h01D6] <= 32'h00300693;
    mem['h01D7] <= 32'hFEC42783;
    mem['h01D8] <= 32'h40F687B3;
    mem['h01D9] <= 32'h00379793;
    mem['h01DA] <= 32'h00F756B3;
    mem['h01DB] <= 32'hFEC42783;
    mem['h01DC] <= 32'hFD842703;
    mem['h01DD] <= 32'h00F707B3;
    mem['h01DE] <= 32'h0FF6F713;
    mem['h01DF] <= 32'h00E78023;
    mem['h01E0] <= 32'hFDC42783;
    mem['h01E1] <= 32'h0547A703;
    mem['h01E2] <= 32'h00300693;
    mem['h01E3] <= 32'hFEC42783;
    mem['h01E4] <= 32'h40F687B3;
    mem['h01E5] <= 32'h00379793;
    mem['h01E6] <= 32'h00F756B3;
    mem['h01E7] <= 32'hFEC42783;
    mem['h01E8] <= 32'h00478793;
    mem['h01E9] <= 32'hFD842703;
    mem['h01EA] <= 32'h00F707B3;
    mem['h01EB] <= 32'h0FF6F713;
    mem['h01EC] <= 32'h00E78023;
    mem['h01ED] <= 32'hFDC42783;
    mem['h01EE] <= 32'h0587A703;
    mem['h01EF] <= 32'h00300693;
    mem['h01F0] <= 32'hFEC42783;
    mem['h01F1] <= 32'h40F687B3;
    mem['h01F2] <= 32'h00379793;
    mem['h01F3] <= 32'h00F756B3;
    mem['h01F4] <= 32'hFEC42783;
    mem['h01F5] <= 32'h00878793;
    mem['h01F6] <= 32'hFD842703;
    mem['h01F7] <= 32'h00F707B3;
    mem['h01F8] <= 32'h0FF6F713;
    mem['h01F9] <= 32'h00E78023;
    mem['h01FA] <= 32'hFDC42783;
    mem['h01FB] <= 32'h05C7A703;
    mem['h01FC] <= 32'h00300693;
    mem['h01FD] <= 32'hFEC42783;
    mem['h01FE] <= 32'h40F687B3;
    mem['h01FF] <= 32'h00379793;
    mem['h0200] <= 32'h00F756B3;
    mem['h0201] <= 32'hFEC42783;
    mem['h0202] <= 32'h00C78793;
    mem['h0203] <= 32'hFD842703;
    mem['h0204] <= 32'h00F707B3;
    mem['h0205] <= 32'h0FF6F713;
    mem['h0206] <= 32'h00E78023;
    mem['h0207] <= 32'hFDC42783;
    mem['h0208] <= 32'h0607A703;
    mem['h0209] <= 32'h00300693;
    mem['h020A] <= 32'hFEC42783;
    mem['h020B] <= 32'h40F687B3;
    mem['h020C] <= 32'h00379793;
    mem['h020D] <= 32'h00F756B3;
    mem['h020E] <= 32'hFEC42783;
    mem['h020F] <= 32'h01078793;
    mem['h0210] <= 32'hFD842703;
    mem['h0211] <= 32'h00F707B3;
    mem['h0212] <= 32'h0FF6F713;
    mem['h0213] <= 32'h00E78023;
    mem['h0214] <= 32'hFDC42783;
    mem['h0215] <= 32'h0647A703;
    mem['h0216] <= 32'h00300693;
    mem['h0217] <= 32'hFEC42783;
    mem['h0218] <= 32'h40F687B3;
    mem['h0219] <= 32'h00379793;
    mem['h021A] <= 32'h00F756B3;
    mem['h021B] <= 32'hFEC42783;
    mem['h021C] <= 32'h01478793;
    mem['h021D] <= 32'hFD842703;
    mem['h021E] <= 32'h00F707B3;
    mem['h021F] <= 32'h0FF6F713;
    mem['h0220] <= 32'h00E78023;
    mem['h0221] <= 32'hFDC42783;
    mem['h0222] <= 32'h0687A703;
    mem['h0223] <= 32'h00300693;
    mem['h0224] <= 32'hFEC42783;
    mem['h0225] <= 32'h40F687B3;
    mem['h0226] <= 32'h00379793;
    mem['h0227] <= 32'h00F756B3;
    mem['h0228] <= 32'hFEC42783;
    mem['h0229] <= 32'h01878793;
    mem['h022A] <= 32'hFD842703;
    mem['h022B] <= 32'h00F707B3;
    mem['h022C] <= 32'h0FF6F713;
    mem['h022D] <= 32'h00E78023;
    mem['h022E] <= 32'hFDC42783;
    mem['h022F] <= 32'h06C7A703;
    mem['h0230] <= 32'h00300693;
    mem['h0231] <= 32'hFEC42783;
    mem['h0232] <= 32'h40F687B3;
    mem['h0233] <= 32'h00379793;
    mem['h0234] <= 32'h00F756B3;
    mem['h0235] <= 32'hFEC42783;
    mem['h0236] <= 32'h01C78793;
    mem['h0237] <= 32'hFD842703;
    mem['h0238] <= 32'h00F707B3;
    mem['h0239] <= 32'h0FF6F713;
    mem['h023A] <= 32'h00E78023;
    mem['h023B] <= 32'hFEC42783;
    mem['h023C] <= 32'h00178793;
    mem['h023D] <= 32'hFEF42623;
    mem['h023E] <= 32'hFEC42703;
    mem['h023F] <= 32'h00300793;
    mem['h0240] <= 32'hE4E7D8E3;
    mem['h0241] <= 32'h00000013;
    mem['h0242] <= 32'h00000013;
    mem['h0243] <= 32'h02C12083;
    mem['h0244] <= 32'h02812403;
    mem['h0245] <= 32'h03010113;
    mem['h0246] <= 32'h00008067;
    mem['h0247] <= 32'hF4010113;
    mem['h0248] <= 32'h0A112E23;
    mem['h0249] <= 32'h0A812C23;
    mem['h024A] <= 32'h0C010413;
    mem['h024B] <= 32'hF4A42623;
    mem['h024C] <= 32'hF4B42423;
    mem['h024D] <= 32'hF4C42223;
    mem['h024E] <= 32'hF7C40793;
    mem['h024F] <= 32'h00078513;
    mem['h0250] <= 32'hA49FF0EF;
    mem['h0251] <= 32'hF7C40793;
    mem['h0252] <= 32'hF4842603;
    mem['h0253] <= 32'hF4C42583;
    mem['h0254] <= 32'h00078513;
    mem['h0255] <= 32'hAB5FF0EF;
    mem['h0256] <= 32'hF5C40713;
    mem['h0257] <= 32'hF7C40793;
    mem['h0258] <= 32'h00070593;
    mem['h0259] <= 32'h00078513;
    mem['h025A] <= 32'hBA1FF0EF;
    mem['h025B] <= 32'hFE042623;
    mem['h025C] <= 32'h0680006F;
    mem['h025D] <= 32'hFEC42783;
    mem['h025E] <= 32'hFF078793;
    mem['h025F] <= 32'h008787B3;
    mem['h0260] <= 32'hF6C7C783;
    mem['h0261] <= 32'hF5840713;
    mem['h0262] <= 32'h00070593;
    mem['h0263] <= 32'h00078513;
    mem['h0264] <= 32'hFA8FF0EF;
    mem['h0265] <= 32'hFEC42783;
    mem['h0266] <= 32'h00179793;
    mem['h0267] <= 32'h00078713;
    mem['h0268] <= 32'hF4442783;
    mem['h0269] <= 32'h00E787B3;
    mem['h026A] <= 32'hF5844703;
    mem['h026B] <= 32'h00E78023;
    mem['h026C] <= 32'hFEC42783;
    mem['h026D] <= 32'h00179793;
    mem['h026E] <= 32'h00178793;
    mem['h026F] <= 32'hF4442703;
    mem['h0270] <= 32'h00F707B3;
    mem['h0271] <= 32'hF5944703;
    mem['h0272] <= 32'h00E78023;
    mem['h0273] <= 32'hFEC42783;
    mem['h0274] <= 32'h00178793;
    mem['h0275] <= 32'hFEF42623;
    mem['h0276] <= 32'hFEC42703;
    mem['h0277] <= 32'h01F00793;
    mem['h0278] <= 32'hF8E7DAE3;
    mem['h0279] <= 32'hF4442783;
    mem['h027A] <= 32'h04078793;
    mem['h027B] <= 32'h00078023;
    mem['h027C] <= 32'h00000013;
    mem['h027D] <= 32'h0BC12083;
    mem['h027E] <= 32'h0B812403;
    mem['h027F] <= 32'h0C010113;
    mem['h0280] <= 32'h00008067;
    mem['h0281] <= 32'h6C6C6548;
    mem['h0282] <= 32'h57202C6F;
    mem['h0283] <= 32'h646C726F;
    mem['h0284] <= 32'h00000021;
    mem['h0285] <= 32'h33323130;
    mem['h0286] <= 32'h37363534;
    mem['h0287] <= 32'h62613938;
    mem['h0288] <= 32'h66656463;
    mem['h0289] <= 32'h00000000;

  end

  always @(posedge clk) mem_data <= mem[mem_addr];

  // ============================================================================

  reg o_ready;

  always @(posedge clk or negedge rstn)
    if (!rstn) o_ready <= 1'd0;
    else o_ready <= valid && ((addr & MEM_ADDR_MASK) != 0);

  // Output connectins
  assign ready    = o_ready;
  assign rdata    = mem_data;
  assign mem_addr = addr[MEM_SIZE_BITS+1:2];

endmodule
